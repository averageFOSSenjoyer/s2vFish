module sKey
(
    input logic [127:0] m,
    output logic [31:0] s0, s1
);

    always_comb begin
        s0[7:0]   = 8'h01 * m[7:0] + 8'hA4 * m[15:8] + 8'h55 * m[23:16] + 8'h87 * m[31:24] + 8'h5A * m[39:32] + 8'h58 * m[47:40] + 8'hDB * m[55:48] + 8'h9E * m[63:56];
        s0[15:8]  = 8'hA4 * m[7:0] + 8'h56 * m[15:8] + 8'h82 * m[23:16] + 8'hF3 * m[31:24] + 8'h1E * m[39:32] + 8'hC6 * m[47:40] + 8'h68 * m[55:48] + 8'hE5 * m[63:56];
        s0[23:16] = 8'h02 * m[7:0] + 8'hA1 * m[15:8] + 8'hFC * m[23:16] + 8'hC1 * m[31:24] + 8'h47 * m[39:32] + 8'hAE * m[47:40] + 8'h3D * m[55:48] + 8'h19 * m[63:56];
        s0[31:24] = 8'hA4 * m[7:0] + 8'h55 * m[15:8] + 8'h87 * m[23:16] + 8'h5A * m[31:24] + 8'h58 * m[39:32] + 8'hDB * m[47:40] + 8'h9E * m[55:48] + 8'h03 * m[63:56];

        s1[7:0]   = 8'h01 * m[71:64] + 8'hA4 * m[79:72] + 8'h55 * m[87:80] + 8'h87 * m[95:88] + 8'h5A * m[103:96] + 8'h58 * m[111:104] + 8'hDB * m[119:112] + 8'h9E * m[127:120];
        s1[15:8]  = 8'hA4 * m[71:64] + 8'h56 * m[79:72] + 8'h82 * m[87:80] + 8'hF3 * m[95:88] + 8'h1E * m[103:96] + 8'hC6 * m[111:104] + 8'h68 * m[119:112] + 8'hE5 * m[127:120];
        s1[23:16] = 8'h02 * m[71:64] + 8'hA1 * m[79:72] + 8'hFC * m[87:80] + 8'hC1 * m[95:88] + 8'h47 * m[103:96] + 8'hAE * m[111:104] + 8'h3D * m[119:112] + 8'h19 * m[127:120];
        s1[31:24] = 8'hA4 * m[71:64] + 8'h55 * m[79:72] + 8'h87 * m[87:80] + 8'h5A * m[95:88] + 8'h58 * m[103:96] + 8'hDB * m[111:104] + 8'h9E * m[119:112] + 8'h03 * m[127:120];
    end

endmodule
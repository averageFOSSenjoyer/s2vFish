// NIOSsoc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module NIOSsoc (
		output wire [31:0] block0_export,    //     block0.export
		output wire [31:0] block1_export,    //     block1.export
		output wire [31:0] block2_export,    //     block2.export
		output wire [31:0] block3_export,    //     block3.export
		input  wire        busy_export,      //       busy.export
		input  wire        clk_clk,          //        clk.clk
		output wire        ende_export,      //       ende.export
		output wire [31:0] key0_export,      //       key0.export
		output wire [31:0] key1_export,      //       key1.export
		output wire [31:0] key2_export,      //       key2.export
		output wire [31:0] key3_export,      //       key3.export
		input  wire [31:0] out0_export,      //       out0.export
		input  wire [31:0] out1_export,      //       out1.export
		input  wire [31:0] out2_export,      //       out2.export
		input  wire [31:0] out3_export,      //       out3.export
		input  wire        reset_reset_n,    //      reset.reset_n
		output wire        reset_1_export,   //    reset_1.export
		output wire        sdram_clk_clk,    //  sdram_clk.clk
		output wire [12:0] sdram_wire_addr,  // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,    //           .ba
		output wire        sdram_wire_cas_n, //           .cas_n
		output wire        sdram_wire_cke,   //           .cke
		output wire        sdram_wire_cs_n,  //           .cs_n
		inout  wire [15:0] sdram_wire_dq,    //           .dq
		output wire [1:0]  sdram_wire_dqm,   //           .dqm
		output wire        sdram_wire_ras_n, //           .ras_n
		output wire        sdram_wire_we_n,  //           .we_n
		output wire        start_export      //      start.export
	);

	wire         sdram_pll_c0_clk;                                            // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_001:clk, sdram:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;              // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;               // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                  // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                 // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;             // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_block0_s1_chipselect;                      // mm_interconnect_0:block0_s1_chipselect -> block0:chipselect
	wire  [31:0] mm_interconnect_0_block0_s1_readdata;                        // block0:readdata -> mm_interconnect_0:block0_s1_readdata
	wire   [1:0] mm_interconnect_0_block0_s1_address;                         // mm_interconnect_0:block0_s1_address -> block0:address
	wire         mm_interconnect_0_block0_s1_write;                           // mm_interconnect_0:block0_s1_write -> block0:write_n
	wire  [31:0] mm_interconnect_0_block0_s1_writedata;                       // mm_interconnect_0:block0_s1_writedata -> block0:writedata
	wire         mm_interconnect_0_block1_s1_chipselect;                      // mm_interconnect_0:block1_s1_chipselect -> block1:chipselect
	wire  [31:0] mm_interconnect_0_block1_s1_readdata;                        // block1:readdata -> mm_interconnect_0:block1_s1_readdata
	wire   [1:0] mm_interconnect_0_block1_s1_address;                         // mm_interconnect_0:block1_s1_address -> block1:address
	wire         mm_interconnect_0_block1_s1_write;                           // mm_interconnect_0:block1_s1_write -> block1:write_n
	wire  [31:0] mm_interconnect_0_block1_s1_writedata;                       // mm_interconnect_0:block1_s1_writedata -> block1:writedata
	wire         mm_interconnect_0_block2_s1_chipselect;                      // mm_interconnect_0:block2_s1_chipselect -> block2:chipselect
	wire  [31:0] mm_interconnect_0_block2_s1_readdata;                        // block2:readdata -> mm_interconnect_0:block2_s1_readdata
	wire   [1:0] mm_interconnect_0_block2_s1_address;                         // mm_interconnect_0:block2_s1_address -> block2:address
	wire         mm_interconnect_0_block2_s1_write;                           // mm_interconnect_0:block2_s1_write -> block2:write_n
	wire  [31:0] mm_interconnect_0_block2_s1_writedata;                       // mm_interconnect_0:block2_s1_writedata -> block2:writedata
	wire         mm_interconnect_0_block3_s1_chipselect;                      // mm_interconnect_0:block3_s1_chipselect -> block3:chipselect
	wire  [31:0] mm_interconnect_0_block3_s1_readdata;                        // block3:readdata -> mm_interconnect_0:block3_s1_readdata
	wire   [1:0] mm_interconnect_0_block3_s1_address;                         // mm_interconnect_0:block3_s1_address -> block3:address
	wire         mm_interconnect_0_block3_s1_write;                           // mm_interconnect_0:block3_s1_write -> block3:write_n
	wire  [31:0] mm_interconnect_0_block3_s1_writedata;                       // mm_interconnect_0:block3_s1_writedata -> block3:writedata
	wire         mm_interconnect_0_key0_s1_chipselect;                        // mm_interconnect_0:key0_s1_chipselect -> key0:chipselect
	wire  [31:0] mm_interconnect_0_key0_s1_readdata;                          // key0:readdata -> mm_interconnect_0:key0_s1_readdata
	wire   [1:0] mm_interconnect_0_key0_s1_address;                           // mm_interconnect_0:key0_s1_address -> key0:address
	wire         mm_interconnect_0_key0_s1_write;                             // mm_interconnect_0:key0_s1_write -> key0:write_n
	wire  [31:0] mm_interconnect_0_key0_s1_writedata;                         // mm_interconnect_0:key0_s1_writedata -> key0:writedata
	wire         mm_interconnect_0_key1_s1_chipselect;                        // mm_interconnect_0:key1_s1_chipselect -> key1:chipselect
	wire  [31:0] mm_interconnect_0_key1_s1_readdata;                          // key1:readdata -> mm_interconnect_0:key1_s1_readdata
	wire   [1:0] mm_interconnect_0_key1_s1_address;                           // mm_interconnect_0:key1_s1_address -> key1:address
	wire         mm_interconnect_0_key1_s1_write;                             // mm_interconnect_0:key1_s1_write -> key1:write_n
	wire  [31:0] mm_interconnect_0_key1_s1_writedata;                         // mm_interconnect_0:key1_s1_writedata -> key1:writedata
	wire         mm_interconnect_0_key2_s1_chipselect;                        // mm_interconnect_0:key2_s1_chipselect -> key2:chipselect
	wire  [31:0] mm_interconnect_0_key2_s1_readdata;                          // key2:readdata -> mm_interconnect_0:key2_s1_readdata
	wire   [1:0] mm_interconnect_0_key2_s1_address;                           // mm_interconnect_0:key2_s1_address -> key2:address
	wire         mm_interconnect_0_key2_s1_write;                             // mm_interconnect_0:key2_s1_write -> key2:write_n
	wire  [31:0] mm_interconnect_0_key2_s1_writedata;                         // mm_interconnect_0:key2_s1_writedata -> key2:writedata
	wire         mm_interconnect_0_key3_s1_chipselect;                        // mm_interconnect_0:key3_s1_chipselect -> key3:chipselect
	wire  [31:0] mm_interconnect_0_key3_s1_readdata;                          // key3:readdata -> mm_interconnect_0:key3_s1_readdata
	wire   [1:0] mm_interconnect_0_key3_s1_address;                           // mm_interconnect_0:key3_s1_address -> key3:address
	wire         mm_interconnect_0_key3_s1_write;                             // mm_interconnect_0:key3_s1_write -> key3:write_n
	wire  [31:0] mm_interconnect_0_key3_s1_writedata;                         // mm_interconnect_0:key3_s1_writedata -> key3:writedata
	wire  [31:0] mm_interconnect_0_out0_s1_readdata;                          // out0:readdata -> mm_interconnect_0:out0_s1_readdata
	wire   [1:0] mm_interconnect_0_out0_s1_address;                           // mm_interconnect_0:out0_s1_address -> out0:address
	wire  [31:0] mm_interconnect_0_out1_s1_readdata;                          // out1:readdata -> mm_interconnect_0:out1_s1_readdata
	wire   [1:0] mm_interconnect_0_out1_s1_address;                           // mm_interconnect_0:out1_s1_address -> out1:address
	wire  [31:0] mm_interconnect_0_out2_s1_readdata;                          // out2:readdata -> mm_interconnect_0:out2_s1_readdata
	wire   [1:0] mm_interconnect_0_out2_s1_address;                           // mm_interconnect_0:out2_s1_address -> out2:address
	wire  [31:0] mm_interconnect_0_out3_s1_readdata;                          // out3:readdata -> mm_interconnect_0:out3_s1_readdata
	wire   [1:0] mm_interconnect_0_out3_s1_address;                           // mm_interconnect_0:out3_s1_address -> out3:address
	wire         mm_interconnect_0_start_s1_chipselect;                       // mm_interconnect_0:start_s1_chipselect -> start:chipselect
	wire  [31:0] mm_interconnect_0_start_s1_readdata;                         // start:readdata -> mm_interconnect_0:start_s1_readdata
	wire   [1:0] mm_interconnect_0_start_s1_address;                          // mm_interconnect_0:start_s1_address -> start:address
	wire         mm_interconnect_0_start_s1_write;                            // mm_interconnect_0:start_s1_write -> start:write_n
	wire  [31:0] mm_interconnect_0_start_s1_writedata;                        // mm_interconnect_0:start_s1_writedata -> start:writedata
	wire         mm_interconnect_0_ende_s1_chipselect;                        // mm_interconnect_0:ende_s1_chipselect -> ende:chipselect
	wire  [31:0] mm_interconnect_0_ende_s1_readdata;                          // ende:readdata -> mm_interconnect_0:ende_s1_readdata
	wire   [1:0] mm_interconnect_0_ende_s1_address;                           // mm_interconnect_0:ende_s1_address -> ende:address
	wire         mm_interconnect_0_ende_s1_write;                             // mm_interconnect_0:ende_s1_write -> ende:write_n
	wire  [31:0] mm_interconnect_0_ende_s1_writedata;                         // mm_interconnect_0:ende_s1_writedata -> ende:writedata
	wire         mm_interconnect_0_reset_s1_chipselect;                       // mm_interconnect_0:reset_s1_chipselect -> reset:chipselect
	wire  [31:0] mm_interconnect_0_reset_s1_readdata;                         // reset:readdata -> mm_interconnect_0:reset_s1_readdata
	wire   [1:0] mm_interconnect_0_reset_s1_address;                          // mm_interconnect_0:reset_s1_address -> reset:address
	wire         mm_interconnect_0_reset_s1_write;                            // mm_interconnect_0:reset_s1_write -> reset:write_n
	wire  [31:0] mm_interconnect_0_reset_s1_writedata;                        // mm_interconnect_0:reset_s1_writedata -> reset:writedata
	wire  [31:0] mm_interconnect_0_busy_s1_readdata;                          // busy:readdata -> mm_interconnect_0:busy_s1_readdata
	wire   [1:0] mm_interconnect_0_busy_s1_address;                           // mm_interconnect_0:busy_s1_address -> busy:address
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [block0:reset_n, block1:reset_n, block2:reset_n, block3:reset_n, busy:reset_n, ende:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, key0:reset_n, key1:reset_n, key2:reset_n, key3:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, out0:reset_n, out1:reset_n, out2:reset_n, out3:reset_n, reset:reset_n, rst_translator:in_reset, sdram_pll:reset, start:reset_n, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	NIOSsoc_block0 block0 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_block0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_block0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_block0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_block0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_block0_s1_readdata),   //                    .readdata
		.out_port   (block0_export)                           // external_connection.export
	);

	NIOSsoc_block0 block1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_block1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_block1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_block1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_block1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_block1_s1_readdata),   //                    .readdata
		.out_port   (block1_export)                           // external_connection.export
	);

	NIOSsoc_block0 block2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_block2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_block2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_block2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_block2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_block2_s1_readdata),   //                    .readdata
		.out_port   (block2_export)                           // external_connection.export
	);

	NIOSsoc_block0 block3 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_block3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_block3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_block3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_block3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_block3_s1_readdata),   //                    .readdata
		.out_port   (block3_export)                           // external_connection.export
	);

	NIOSsoc_busy busy (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_busy_s1_readdata), //                    .readdata
		.in_port  (busy_export)                         // external_connection.export
	);

	NIOSsoc_ende ende (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ende_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ende_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ende_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ende_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ende_s1_readdata),   //                    .readdata
		.out_port   (ende_export)                           // external_connection.export
	);

	NIOSsoc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	NIOSsoc_block0 key0 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_key0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key0_s1_readdata),   //                    .readdata
		.out_port   (key0_export)                           // external_connection.export
	);

	NIOSsoc_block0 key1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_key1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key1_s1_readdata),   //                    .readdata
		.out_port   (key1_export)                           // external_connection.export
	);

	NIOSsoc_block0 key2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_key2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key2_s1_readdata),   //                    .readdata
		.out_port   (key2_export)                           // external_connection.export
	);

	NIOSsoc_block0 key3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_key3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key3_s1_readdata),   //                    .readdata
		.out_port   (key3_export)                           // external_connection.export
	);

	NIOSsoc_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	NIOSsoc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	NIOSsoc_out0 out0 (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_out0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_out0_s1_readdata), //                    .readdata
		.in_port  (out0_export)                         // external_connection.export
	);

	NIOSsoc_out0 out1 (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_out1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_out1_s1_readdata), //                    .readdata
		.in_port  (out1_export)                         // external_connection.export
	);

	NIOSsoc_out0 out2 (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_out2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_out2_s1_readdata), //                    .readdata
		.in_port  (out2_export)                         // external_connection.export
	);

	NIOSsoc_out0 out3 (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_out3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_out3_s1_readdata), //                    .readdata
		.in_port  (out3_export)                         // external_connection.export
	);

	NIOSsoc_ende reset (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reset_s1_readdata),   //                    .readdata
		.out_port   (reset_1_export)                         // external_connection.export
	);

	NIOSsoc_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	NIOSsoc_sdram_pll sdram_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                   //                    c1.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.c2                 (),                                                //           (terminated)
		.c3                 (),                                                //           (terminated)
		.c4                 (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (3'b000),                                          //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	NIOSsoc_ende start (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_s1_readdata),   //                    .readdata
		.out_port   (start_export)                           // external_connection.export
	);

	NIOSsoc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	NIOSsoc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                            //                             sdram_pll_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                          //        sdram_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.block0_s1_address                              (mm_interconnect_0_block0_s1_address),                         //                                block0_s1.address
		.block0_s1_write                                (mm_interconnect_0_block0_s1_write),                           //                                         .write
		.block0_s1_readdata                             (mm_interconnect_0_block0_s1_readdata),                        //                                         .readdata
		.block0_s1_writedata                            (mm_interconnect_0_block0_s1_writedata),                       //                                         .writedata
		.block0_s1_chipselect                           (mm_interconnect_0_block0_s1_chipselect),                      //                                         .chipselect
		.block1_s1_address                              (mm_interconnect_0_block1_s1_address),                         //                                block1_s1.address
		.block1_s1_write                                (mm_interconnect_0_block1_s1_write),                           //                                         .write
		.block1_s1_readdata                             (mm_interconnect_0_block1_s1_readdata),                        //                                         .readdata
		.block1_s1_writedata                            (mm_interconnect_0_block1_s1_writedata),                       //                                         .writedata
		.block1_s1_chipselect                           (mm_interconnect_0_block1_s1_chipselect),                      //                                         .chipselect
		.block2_s1_address                              (mm_interconnect_0_block2_s1_address),                         //                                block2_s1.address
		.block2_s1_write                                (mm_interconnect_0_block2_s1_write),                           //                                         .write
		.block2_s1_readdata                             (mm_interconnect_0_block2_s1_readdata),                        //                                         .readdata
		.block2_s1_writedata                            (mm_interconnect_0_block2_s1_writedata),                       //                                         .writedata
		.block2_s1_chipselect                           (mm_interconnect_0_block2_s1_chipselect),                      //                                         .chipselect
		.block3_s1_address                              (mm_interconnect_0_block3_s1_address),                         //                                block3_s1.address
		.block3_s1_write                                (mm_interconnect_0_block3_s1_write),                           //                                         .write
		.block3_s1_readdata                             (mm_interconnect_0_block3_s1_readdata),                        //                                         .readdata
		.block3_s1_writedata                            (mm_interconnect_0_block3_s1_writedata),                       //                                         .writedata
		.block3_s1_chipselect                           (mm_interconnect_0_block3_s1_chipselect),                      //                                         .chipselect
		.busy_s1_address                                (mm_interconnect_0_busy_s1_address),                           //                                  busy_s1.address
		.busy_s1_readdata                               (mm_interconnect_0_busy_s1_readdata),                          //                                         .readdata
		.ende_s1_address                                (mm_interconnect_0_ende_s1_address),                           //                                  ende_s1.address
		.ende_s1_write                                  (mm_interconnect_0_ende_s1_write),                             //                                         .write
		.ende_s1_readdata                               (mm_interconnect_0_ende_s1_readdata),                          //                                         .readdata
		.ende_s1_writedata                              (mm_interconnect_0_ende_s1_writedata),                         //                                         .writedata
		.ende_s1_chipselect                             (mm_interconnect_0_ende_s1_chipselect),                        //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.key0_s1_address                                (mm_interconnect_0_key0_s1_address),                           //                                  key0_s1.address
		.key0_s1_write                                  (mm_interconnect_0_key0_s1_write),                             //                                         .write
		.key0_s1_readdata                               (mm_interconnect_0_key0_s1_readdata),                          //                                         .readdata
		.key0_s1_writedata                              (mm_interconnect_0_key0_s1_writedata),                         //                                         .writedata
		.key0_s1_chipselect                             (mm_interconnect_0_key0_s1_chipselect),                        //                                         .chipselect
		.key1_s1_address                                (mm_interconnect_0_key1_s1_address),                           //                                  key1_s1.address
		.key1_s1_write                                  (mm_interconnect_0_key1_s1_write),                             //                                         .write
		.key1_s1_readdata                               (mm_interconnect_0_key1_s1_readdata),                          //                                         .readdata
		.key1_s1_writedata                              (mm_interconnect_0_key1_s1_writedata),                         //                                         .writedata
		.key1_s1_chipselect                             (mm_interconnect_0_key1_s1_chipselect),                        //                                         .chipselect
		.key2_s1_address                                (mm_interconnect_0_key2_s1_address),                           //                                  key2_s1.address
		.key2_s1_write                                  (mm_interconnect_0_key2_s1_write),                             //                                         .write
		.key2_s1_readdata                               (mm_interconnect_0_key2_s1_readdata),                          //                                         .readdata
		.key2_s1_writedata                              (mm_interconnect_0_key2_s1_writedata),                         //                                         .writedata
		.key2_s1_chipselect                             (mm_interconnect_0_key2_s1_chipselect),                        //                                         .chipselect
		.key3_s1_address                                (mm_interconnect_0_key3_s1_address),                           //                                  key3_s1.address
		.key3_s1_write                                  (mm_interconnect_0_key3_s1_write),                             //                                         .write
		.key3_s1_readdata                               (mm_interconnect_0_key3_s1_readdata),                          //                                         .readdata
		.key3_s1_writedata                              (mm_interconnect_0_key3_s1_writedata),                         //                                         .writedata
		.key3_s1_chipselect                             (mm_interconnect_0_key3_s1_chipselect),                        //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.out0_s1_address                                (mm_interconnect_0_out0_s1_address),                           //                                  out0_s1.address
		.out0_s1_readdata                               (mm_interconnect_0_out0_s1_readdata),                          //                                         .readdata
		.out1_s1_address                                (mm_interconnect_0_out1_s1_address),                           //                                  out1_s1.address
		.out1_s1_readdata                               (mm_interconnect_0_out1_s1_readdata),                          //                                         .readdata
		.out2_s1_address                                (mm_interconnect_0_out2_s1_address),                           //                                  out2_s1.address
		.out2_s1_readdata                               (mm_interconnect_0_out2_s1_readdata),                          //                                         .readdata
		.out3_s1_address                                (mm_interconnect_0_out3_s1_address),                           //                                  out3_s1.address
		.out3_s1_readdata                               (mm_interconnect_0_out3_s1_readdata),                          //                                         .readdata
		.reset_s1_address                               (mm_interconnect_0_reset_s1_address),                          //                                 reset_s1.address
		.reset_s1_write                                 (mm_interconnect_0_reset_s1_write),                            //                                         .write
		.reset_s1_readdata                              (mm_interconnect_0_reset_s1_readdata),                         //                                         .readdata
		.reset_s1_writedata                             (mm_interconnect_0_reset_s1_writedata),                        //                                         .writedata
		.reset_s1_chipselect                            (mm_interconnect_0_reset_s1_chipselect),                       //                                         .chipselect
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),               //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),                 //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),                  //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),              //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata),             //                                         .writedata
		.start_s1_address                               (mm_interconnect_0_start_s1_address),                          //                                 start_s1.address
		.start_s1_write                                 (mm_interconnect_0_start_s1_write),                            //                                         .write
		.start_s1_readdata                              (mm_interconnect_0_start_s1_readdata),                         //                                         .readdata
		.start_s1_writedata                             (mm_interconnect_0_start_s1_writedata),                        //                                         .writedata
		.start_s1_chipselect                            (mm_interconnect_0_start_s1_chipselect),                       //                                         .chipselect
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)        //                                         .readdata
	);

	NIOSsoc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (sdram_pll_c0_clk),                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
